`ifndef __FREE_LIST_V__
`define __FREE_LIST_V__

`define BIN_LEN 6
`define OUT_BIN_LEN 6
`define SC_LEN 64
`define BIN_WIDTH 3


`define KERNEL_WIDTH 2
`define KERNEL_HEIGHT 2
`define INPUT_WIDTH 4
`define INPUT_HEIGHT 4
`define INPUT_WIDTH_LOG 2
`define INPUT_HEIGHT_LOG 2

`endif
